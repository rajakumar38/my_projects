//class 
//class is a user defined data type that contains data members and methods
//class are dynamically allocated and destroyed
//properties and methods are accesed after creating an object.
//accesed by using handle
//sv supports nested classes
