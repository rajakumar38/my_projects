/*

this is uma

*/



module top;

initial begin


$display("=================this is uma===============================:");

end

endmodule
